--! \addtogroup PropHeatFsm2x1Mode_Module
--! @{
--! \addtogroup PropHeatFsm2x1Mode_Result
--! @{
--! @brief Testbench for the PropHeatFsm2x1Mode module
--! @page PropHeatFsm2x1Mode
--! @section PropHeatFsm2x1Mode Result of tests
--! <b>State machine test - Full run. Test Name: state_machine_full_en3_tb</b> \n
--! EN3 and RstTmr_TB shall be high(1) and low(0) according to the steps defined in HHLR_452. \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_452 |
--! | Tests HHLR_453 |
--! | Tests DHHLR_460 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.state_machine_full_en3_tb_1.png state_machine_full_en3_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.state_machine_full_en3_tb_1.png state_machine_full_en3_tb_1 width=16cm
--! \n
--! State machine test - State 0 - EN1_TB, EN2_TB, EN3_TB and EN4_TB were low(0) and RstTmr_TB was high(1): \b PASS \n \n
--! State machine test - State 1 - EN2_TB was low(0) and RstTmr_TB was low(0): \b PASS \n \n
--! State machine test - State 2 - EN2_TB was high(1) and RstTmr_TB was high(1): \b PASS \n \n
--! State machine test - State 3 - EN3_TB was low(0) and RstTmr_TB was low(0): \b PASS \n \n
--! State machine test - State 4 - EN3_TB was high(1) and RstTmr_TB was high(1): \b PASS \n \n
--! State machine test - State 1 - EN3_TB was low(0) and RstTmr_TB was low(0): \b PASS \n \n
--! <b>Self test override channel one active. Test Name: self_test_overr_ch1_tb</b> \n
--! SelfTestOverrideCh1_TB shall enable EN1_TB regardless of other input states. \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_454 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch1_tb_1.png self_test_overr_ch1_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch1_tb_1.png self_test_overr_ch1_tb_1 width=16cm
--! \n
--! EN1_TB was set to high(1) by SelfTestOverrideCh1_TB and remained high(1) while all other inputs where toggled: \b PASS \n \n
--! <b>Self test override channel two active. Test Name: self_test_overr_ch2_tb</b> \n
--! SelfTestOverrideCh2_TB shall enable EN2_TB regardless of other input states. \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_455 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch2_tb_1.png self_test_overr_ch2_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch2_tb_1.png self_test_overr_ch2_tb_1 width=16cm
--! \n
--! EN2_TB was set to high(1) by SelfTestOverrideCh2_TB and remained high(1) while all other inputs where toggled: \b PASS \n \n
--! <b>Self test override channel three active. Test Name: self_test_overr_ch3_tb</b> \n
--! SelfTestOverrideCh3_TB shall enable EN3_TB regardless of other input states. \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_456 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch3_tb_1.png self_test_overr_ch3_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch3_tb_1.png self_test_overr_ch3_tb_1 width=16cm
--! \n
--! EN3_TB was set to high(1) by SelfTestOverrideCh3_TB and remained high(1) while all other inputs where toggled: \b PASS \n \n
--! <b>Self test override channel four active. Test Name: self_test_overr_ch4_tb</b> \n
--! SelfTestOverrideCh4_TB shall enable EN4_TB regardless of other input states. \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_457 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch4_tb_1.png self_test_overr_ch4_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_overr_ch4_tb_1.png self_test_overr_ch4_tb_1 width=16cm
--! \n
--! EN4_TB was set to high(1) by SelfTestOverrideCh4_TB and remained high(1) while all other inputs where toggled: \b PASS \n \n
--! <b>Self test override from state one. Test Name: self_test_override_from_state_one</b> \n
--! SelfTestOverrideCh1_TB, SelfTestOverrideCh2_TB, SelfTestOverrideCh3_TB and SelfTestOverrideCh4_TB are switched to high(1) in state one, the respective output must get active(1). \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_452 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_override_from_state_one_1.png self_test_override_from_state_one_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_override_from_state_one_1.png self_test_override_from_state_one_1 width=16cm
--! \n
--! EN1_TB, EN2_TB, EN3_TB and EN4_TB are active(1): \b PASS \n \n
--! <b>Self test override from state three. Test Name: self_test_override_from_state_three</b> \n
--! SelfTestOverrideCh1_TB, SelfTestOverrideCh2_TB, SelfTestOverrideCh3_TB and SelfTestOverrideCh4_TB are switched to high(1) in state three, the respective output must get active(1). \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_452 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_override_from_state_three_1.png self_test_override_from_state_three_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_override_from_state_three_1.png self_test_override_from_state_three_1 width=16cm
--! \n
--! EN1_TB, EN2_TB, EN3_TB and EN4_TB are active(1): \b PASS \n \n
--! <b>Self test override from state four. Test Name: self_test_override_from_state_four</b> \n
--! SelfTestOverrideCh1_TB, SelfTestOverrideCh2_TB, SelfTestOverrideCh3_TB and SelfTestOverrideCh4_TB are switched to high(1) in state four, the respective output must get active(1). \n
--! \n
--! | Requirement(s) Covered |
--! | :-: |
--! | Tests HHLR_452 |
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.self_test_override_from_state_four_1.png self_test_override_from_state_four_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.self_test_override_from_state_four_1.png self_test_override_from_state_four_1 width=16cm
--! \n
--! EN1_TB, EN2_TB, EN3_TB and EN4_TB are active(1): \b PASS \n \n
--! <b>Transition coverage - state1 to state0 test. Test Name: trans_state1_to_state0_tb</b> \n
--! RstTmr_TB shall change from low(0) in state1 to high(1) in state0. \n
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.trans_state1_to_state0_tb_1.png trans_state1_to_state0_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.trans_state1_to_state0_tb_1.png trans_state1_to_state0_tb_1 width=16cm
--! \n
--! RstTmr_TB changed from state1 low(0) to state0 high(1): \b PASS \n \n
--! <b>Transition coverage - state3 to state0 test. Test Name: trans_state3_to_state0_tb</b> \n
--! RstTmr_TB shall change from low(0) in state3 to high(1) in state0. \n
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.trans_state3_to_state0_tb_1.png trans_state3_to_state0_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.trans_state3_to_state0_tb_1.png trans_state3_to_state0_tb_1 width=16cm
--! \n
--! RstTmr_TB changed from state3 low(0) to state0 high(1): \b PASS \n \n
--! <b>Transition coverage - state4 to state0 test. Test Name: trans_state4_to_state0_tb</b> \n
--! RstTmr_TB shall change from low(0) in state4 to high(1) in state0. \n
--! \n
--! @image html lib.e_propheatfsm2x1modequalification_tb.trans_state4_to_state0_tb_1.png trans_state4_to_state0_tb_1 width=1000
--! @image latex lib.e_propheatfsm2x1modequalification_tb.trans_state4_to_state0_tb_1.png trans_state4_to_state0_tb_1 width=16cm
--! \n
--! RstTmr_TB changed from state4 low(0) to state0 low(0): \b PASS \n \n
--! \n \n
entity e_propheatfsm2x1modeLog is 
end e_propheatfsm2x1modeLog;
architecture a_propheatfsm2x1modeLog of e_propheatfsm2x1modeLog is
begin
end a_propheatfsm2x1modeLog;
--! @}
--! @}
